LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

ENTITY ram_32_64 IS
PORT(
clk:IN STD_LOGIC;
wr:IN STD_LOGIC;
addr_in:IN STD_LOGIC_VECTOR(4 DOWNTO 0);
addr_out:IN STD_LOGIC_VECTOR(4 DOWNTO 0);
ram_in:IN STD_LOGIC_VECTOR(63 DOWNTO 0);
ram_out:OUT STD_LOGIC_VECTOR(63 DOWNTO 0)
);
END ENTITY;

ARCHITECTURE Behavioral OF ram_32_64 IS
SUBTYPE WORD IS STD_LOGIC_VECTOR(63 DOWNTO 0);
TYPE MEMORY IS ARRAY(32 DOWNTO 0) OF WORD;
SIGNAL ram_mem:MEMORY;

BEGIN

PROCESS(clk)
 BEGIN
  IF(clk'EVENT AND clk='1')THEN
    
	  IF(wr='1')THEN
	     ram_mem(CONV_INTEGER(addr_in))<=ram_in;
	  ELSE
	     ram_out<= ram_mem(CONV_INTEGER(addr_out));
	  END IF;
 
  END IF;
END PROCESS;
END Behavioral;
